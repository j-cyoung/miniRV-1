module shift(
        input   wire            dir,    // dir=0 ��ʾ����, dir=1 ��ʾ����
        input   wire            al,     // al=1 ��ʾ��������
        input   wire    [31:0]  a,
        input   wire    [4:0]   b,
        output  reg     [31:0]  c
    );

always@(*) begin
    if (dir)    // ����
        case(b)
            5'd0:   c = a;
            5'd1 :  c = {{ 1{al&a[31]}}, a[31: 1]};
            5'd2 :  c = {{ 2{al&a[31]}}, a[31: 2]};
            5'd3 :  c = {{ 3{al&a[31]}}, a[31: 3]};
            5'd4 :  c = {{ 4{al&a[31]}}, a[31: 4]};
            5'd5 :  c = {{ 5{al&a[31]}}, a[31: 5]};
            5'd6 :  c = {{ 6{al&a[31]}}, a[31: 6]};
            5'd7 :  c = {{ 7{al&a[31]}}, a[31: 7]};
            5'd8 :  c = {{ 8{al&a[31]}}, a[31: 8]};
            5'd9 :  c = {{ 9{al&a[31]}}, a[31: 9]};
            5'd10:  c = {{10{al&a[31]}}, a[31:10]};               
            5'd11:  c = {{11{al&a[31]}}, a[31:11]};
            5'd12:  c = {{12{al&a[31]}}, a[31:12]};
            5'd13:  c = {{13{al&a[31]}}, a[31:13]};
            5'd14:  c = {{14{al&a[31]}}, a[31:14]};
            5'd15:  c = {{15{al&a[31]}}, a[31:15]};
            5'd16:  c = {{16{al&a[31]}}, a[31:16]};
            5'd17:  c = {{17{al&a[31]}}, a[31:17]};
            5'd18:  c = {{18{al&a[31]}}, a[31:18]};
            5'd19:  c = {{19{al&a[31]}}, a[31:19]};
            5'd20:  c = {{20{al&a[31]}}, a[31:20]};
            5'd21:  c = {{21{al&a[31]}}, a[31:21]};
            5'd22:  c = {{22{al&a[31]}}, a[31:22]};
            5'd23:  c = {{23{al&a[31]}}, a[31:23]};
            5'd24:  c = {{24{al&a[31]}}, a[31:24]};
            5'd25:  c = {{25{al&a[31]}}, a[31:25]};
            5'd26:  c = {{26{al&a[31]}}, a[31:26]};
            5'd27:  c = {{27{al&a[31]}}, a[31:27]};
            5'd28:  c = {{28{al&a[31]}}, a[31:28]};
            5'd29:  c = {{29{al&a[31]}}, a[31:29]};
            5'd30:  c = {{30{al&a[31]}}, a[31:30]};
            5'd31:  c = {{31{al&a[31]}}, a[31:31]};
        default:
            c = {32{al&a[31]}};
        endcase
    else    // ����
        case(b)
            5'd0:   c = a;
            5'd1:   c = {a[30: 0], 1'b0};
            5'd2:   c = {a[29: 0], 2'b0};
            5'd3:   c = {a[28: 0], 3'b0};
            5'd4:   c = {a[27: 0], 4'b0};
            5'd5:   c = {a[26: 0], 5'b0};
            5'd6:   c = {a[25: 0], 6'b0};
            5'd7:   c = {a[24: 0], 7'b0};
            5'd8:   c = {a[23: 0], 8'b0};
            5'd9:   c = {a[22: 0], 9'b0};
            5'd10:  c = {a[21: 0],10'b0};               
            5'd11:  c = {a[20: 0],11'b0};
            5'd12:  c = {a[19: 0],12'b0};
            5'd13:  c = {a[18: 0],13'b0};
            5'd14:  c = {a[17: 0],14'b0};
            5'd15:  c = {a[16: 0],15'b0};
            5'd16:  c = {a[15: 0],16'b0};
            5'd17:  c = {a[14: 0],17'b0};
            5'd18:  c = {a[13: 0],18'b0};
            5'd19:  c = {a[12: 0],19'b0};
            5'd20:  c = {a[11: 0],20'b0};
            5'd21:  c = {a[10: 0],21'b0};
            5'd22:  c = {a[ 9: 0],22'b0};
            5'd23:  c = {a[ 8: 0],23'b0};
            5'd24:  c = {a[ 7: 0],24'b0};
            5'd25:  c = {a[ 6: 0],25'b0};
            5'd26:  c = {a[ 5: 0],26'b0};
            5'd27:  c = {a[ 4: 0],27'b0};
            5'd28:  c = {a[ 3: 0],28'b0};
            5'd29:  c = {a[ 2: 0],29'b0};
            5'd30:  c = {a[ 1: 0],30'b0};
            5'd31:  c = {a[ 0: 0],31'b0};
        default:
            c = 32'b0;
        endcase
end
    
endmodule